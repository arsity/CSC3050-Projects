//~ `New testbench
`timescale  1ns / 1ps

module tb_alu;

// alu Parameters
parameter PERIOD  = 10;


// alu Inputs
reg   [31:0]  instruction;
reg   [31:0]  regA;
reg   [31:0]  regB;

// alu Outputs
wire  [31:0]  result;
wire  [2:0]  flags;

alu  u_alu (instruction, regA, regB, result, flags);

initial begin
    $display(" instruction : reg_A : reg_B : result : flags ");
    $monitor(" %h : %h : %h : %h : %b ", instruction, regA, regB, result, flags);


    // add
    #10 instruction   <= 32'b000000_00000_00001_00011_00000_100000    ;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000  ;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000  ;
    
    $display("add");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00011_00000_100000    ;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;

    #10 instruction   <= 32'b000000_00000_00001_00011_00000_100000    ;
    regA              <= 32'b0100_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b0100_0000_0000_0000_0000_0000_0000_0001  ;

    #10 instruction   <= 32'b000000_00000_00001_00011_00000_100000    ;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_1101_1101  ;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_0010_0011  ;

    #10 instruction   <= 32'b000000_00000_00001_00011_00000_100000    ;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0101_1101  ;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_0010_0011  ;


    //addi
    #10 instruction   <= 32'b001000_00000_00001_1000000000100000      ;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;
    
    $display("addi");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b001000_00000_00001_0000000000100010      ;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;

    #10 instruction   <= 32'b001000_00000_00001_0000000000100000      ;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;

    #10 instruction   <= 32'b001000_00000_00001_0000000000100000      ;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0010_0001  ;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;


    //addu
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100001    ;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_1001  ;
    
    $display("addu");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100001    ;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001  ;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100001    ;
    regA              <= 32'b0100_0000_0000_0000_0000_0000_0000_0001  ;
    regB              <= 32'b0100_0000_0000_0000_0000_0000_0000_0001  ;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100001    ;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_1101_1101  ;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_0010_0011  ;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100001    ;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0101_1101  ;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_0010_0011  ;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100001    ;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000  ;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000  ;


    //addiu
    #10 instruction   <= 32'b001001_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("addiu");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b001001_00000_00001_1000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;

    #10 instruction   <= 32'b001001_00000_00001_0000000000000000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;


    //sub
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100010;
    regA              <= 32'b1111_0000_0000_0000_0000_0000_0101_1101;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("sub");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100010;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0111_0000_0000_0000_0000_0000_0101_1101;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100010;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1111_0000_0000_0000_0000_0000_0101_1101;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100010;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;


    //subu
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100011;
    regA              <= 32'b0111_0000_0000_0000_0000_0000_0101_1101;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("subu");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100011;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0111_0000_0000_0000_0000_0000_0101_1101;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100011;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1111_0000_0000_0000_0000_0000_0101_1101;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100011;
    regA              <= 32'b0000_0000_0000_0000_0000_1000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0101_1101;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100011;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;


    //and
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100100;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    
    $display("and");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100100;
    regA              <= 32'b1000_0000_1001_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_1001_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100100;
    regA              <= 32'b1000_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100100;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //andi
    #10 instruction   <= 32'b001100_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("andi");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b001100_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b001100_00000_00001_1000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //nor
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100111;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    
    $display("nor");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100111;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100111;
    regA              <= 32'b1000_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100111;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //or
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_100101;
    regA              <= 32'b1111_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;
    
    $display("or");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_100101;
    regA              <= 32'b0100_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;

    #10 instruction   <= 32'b000000_00000_00001_00001_11000_100101;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;


    //ori
    #10 instruction   <= 32'b001101_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("ori");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b001101_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b001101_00000_00001_0000000000000000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //xor
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100110;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    
    $display("xor");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100110;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100110;
    regA              <= 32'b1000_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_100110;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //xori
    #10 instruction   <= 32'b001110_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("xori");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b001110_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b001110_00000_00001_1000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //beq/bne
    #10 instruction   <= 32'b000100_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("beq/bne");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000100_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b000100_00000_00001_1000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //slt
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101010;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    
    $display("slt");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101010;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101010;
    regA              <= 32'b0100_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101010;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //slti
    #10 instruction   <= 32'b001010_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("slti");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b001010_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b001010_00000_00001_1000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //sltu
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101011;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    
    $display("sltu");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101011;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101011;
    regA              <= 32'b1000_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;

    #10 instruction   <= 32'b000000_00000_00001_00001_00000_101011;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //stliu
    #10 instruction   <= 32'b001011_00000_00001_0000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("stliu");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b001011_00000_00001_0000000000010000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b001011_00000_00001_1000000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b001011_00000_00001_1000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //sw
    #10 instruction   <= 32'b101011_00000_00001_0001000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("sw");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b101011_00000_00001_0000100000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b101011_00000_00001_1000000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //lw
    #10 instruction   <= 32'b100011_00000_00001_0000010000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
    
    $display("lw");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b100011_00000_00001_0001000000100000;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;

    #10 instruction   <= 32'b100011_00000_00001_0010000000100000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;


    //sll
    #10 instruction   <= 32'b000000_00000_00001_00001_00100_000000;
    regA              <= 32'b1111_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;
    $display("sll");
    $display(" instruction : reg_A : reg_B : result : flags ");
    #10 instruction   <= 32'b000000_00000_00001_00001_01000_000000;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //sllv
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_000100;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0010_0010;
    
    $display("sllv");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_000100;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;


    //srl
    #10 instruction   <= 32'b000000_00000_00001_00001_01000_000010;
    regA              <= 32'b1111_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;
    
    $display("srl");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_01000_000010;
    regA              <= 32'b0100_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //srlv
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_000110;
    regA              <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    
    $display("srlv");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_000110;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0000_0110;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;


    //sra
    #10 instruction   <= 32'b000000_00000_00001_00001_01000_000011;
    regA              <= 32'b1111_1100_0010_0000_0000_0000_0000_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0011_0010;
    
    $display("sra");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_01000_000011;
    regA              <= 32'b0100_0000_0000_0000_0000_0000_0000_0000;
    regB              <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;


    //srav
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_000111;
    regA              <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    
    $display("srav");
    $display(" instruction : reg_A : reg_B : result : flags ");
    
    #10 instruction   <= 32'b000000_00000_00001_00001_11000_000111;
    regA              <= 32'b0000_0000_0000_0000_0001_0000_0000_0110;
    regB              <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;

    
    #10 $finish;
end
endmodule